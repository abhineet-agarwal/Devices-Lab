*RN142_RT
.MODEL DRN142S D(IS=127.76E-12 N=1.7346 RS=.1581 IKF=.14089 
+ CJO=385.59E-15 M=.11823 VJ=.78827 ISR=139.38E-12 NR=3 BV=60 TT=275.00E-9)

d1 1 2 DRN142S
r1 2 0 1000
vin 1 0 pulse(0 2 0 1n 1n 0.167u 0.333u)

.tran 0.1n 0.4u                       

.control
run
plot -i(vin) xlimit 0u 0.4u

wrdata diode_recovery.csv time i(vin)
                
.endc

.end