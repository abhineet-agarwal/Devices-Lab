* Solar Cell SPICE Subcircuit Data
.subckt solar_cell PX NX
*IL is photo generated current (keep only 1 of the next 3 lines, whichever is necessary)
*IL NX TMP dc 0e-3
*IL NX TMP dc 8e-3
IL NX TMP dc 10e-3

d1 TMP NX diode
.model diode d (is=(1e-13) n=1)

d2 TMP NX diode2
.model diode2 d (is=(2e-6) n=2)

rs TMP PX 10
rsh TMP NX 1e3

.ends solar_cell

* Main Circuit
* Resistance load connected to the solar cell
r1 2 0 100

* Instantiate the solar cell subcircuit
x1 1 2 solar_cell

* Independent DC source whose voltage is to be varied
vin 1 0 dc 0

* DC Analysis on source vin, to vary from -2 to 2V in 0.01V steps
.dc vin -2 2 0.01

* Control commands for running the simulation
.control
run
* Plot the current through R1 (V(2)/100) vs. the voltage across the solar cell (V(1)-V(2))
plot (v(2)/100) vs v(1)-v(2)
.endc
.end
