*blue_led
.include E:/Devices_Lab/blue_5mm.txt

d1 1 2 BLUE 
r1 2 0 100
vin 1 0 dc
.dc vin 0 5 0.01
.control
run
plot ln(V(2)/100)
.endc
.end